`ifndef ELINK_CONSTANTS_V_
 `define ELINK_CONSTANTS_V_

 `define CFG_TARGET "XILINX"  // default hard macro target
                              // see also "GENERIC", "ALTERA", "ASIC"
 `define CFG_ASIC=0
 `define CFG_PLATFORM=\"ZYNQ\"
`endif
